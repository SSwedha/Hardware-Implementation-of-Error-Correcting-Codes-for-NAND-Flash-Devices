package rm_encoder;
import Vector :: *;
import FIFOF::*;
//(*doc = "note: The architecture is as follows- There is an overall interface "Encoder". It has to sub-interfaces, one to receive input (message) and one to send output (codeword). There is a module to which the interface "encoder" is tied to. Using this module, valid codewords are generated. " *)

//(*doc = "ifc: Overall block of encoder" *)
interface Ifc_rm_encoder;
	//(*doc = "subifc: Subifc_Enc_In takes input(message) from the source "*)
	interface Subifc_Enc_In subifc_in;
	//(*doc = "subifc: Subifc_Enc_Out sends output(codeword) through the channel "*)
	interface Subifc_Enc_Out subifc_out;
endinterface: Ifc_rm_encoder

interface Subifc_Enc_In;
	//(*doc = "method: This Action method receives message(247 bits) from the source "*)
	method Action ma_get_message(Bit#(247) lv_message_in);
endinterface: Subifc_Enc_In

interface Subifc_Enc_Out;
	//(*doc = "method: This ActionValue method sends codeword(256 bits) to the channel "*)
	method ActionValue#(Bit#(256)) mav_tx_codeword;
endinterface: Subifc_Enc_Out

//(*doc = "func:  This function performs matrix multiplication. It multiplies the row vector message to each column of generator matrix. Row vector codeword of 256 bits is returned. " *)
function Bit#(256) fn_mul(Vector#(247,Bit#(256)) v_matrix, Bit#(247) lv_message);
  Bit#(256) lv_codeword = 256'b0;
  //(*doc = "note: The matrix multiplication is from MSB to LSB. Hence the generator matrix can be thought of in this form:)
  
  //(*doc = "note: | g255,0   | g254,0	 | g253,0   |...| g2,0   | g1,0   | g0,0   | "*)
  //(*doc = "note: | g255,1   | g254,1   | g253,1   |...| g2,1   | g1,1   | g0,1   | "*)
  //(*doc = "note: |  .       |  .       |  .       |...|  .     |  .     |  .     | "*)
  //(*doc = "note: |  .       |  .       |  .       |...|  .     |  .     |  .     | "*)
  //(*doc = "note: |  .       |  .       |  .       |...|  .     |  .     |  .     | "*)
  //(*doc = "note: | g255,245 | g254,245 | g253,245 |...| g2,245 | g1,245 | g0,245 | "*)
  //(*doc = "note: | g255,246 | g254,246 | g253,246 |...| g2,246 | g1,246 | g0,246 | "*)
  //(*doc = "note: Thus the coloumn index must start from 255 and decrease till 0. However, the row index can start from 0 or 247. In this case, we are starting from 0. "*)
  for(Integer lv_j=255;lv_j>0;lv_j=lv_j-1)
  begin
  	for(Integer lv_i=0;lv_i<247;lv_i=lv_i+1)
  	begin
  	//(*doc = "note: When an element of column of the matrix is 1, we will XOR the value of 246-i th bit of message vector with the previously stored value of codeword in the jth location. We need to XOR to do mod2 addition. "*)
  		if(v_matrix[lv_i][lv_j] == 1)
  		 //(*doc ="note: We are taking 246-i th bit of message because we need to maintain the order of codeword from MSB to LSB and not the other way around. This can be avoided by making the i loop start from 246 and decreasing it to 0. "*)
  			lv_codeword[lv_j] = lv_codeword[lv_j]^lv_message[246-lv_i];
  	end
  end
  return lv_codeword;
endfunction

(*synthesize*)
(*doc = "module: Encoder module " *)
module mk_rm_encoder (Ifc_rm_encoder);

	(*doc = "fifo:  To store the codeword after the parity bits are generated " *)
	FIFOF#(Bit#(256)) ff_output <- mkFIFOF();
	
	//(*doc = "note:  To store the rows of generator matrix as vector of 247 elements, each with size of 256 bits. " *)
	Vector#(247,Bit#(256)) v_gen;
	
//(*doc = "note: The generator matrix has been generated using the c++ program. "*)
v_gen[0]=256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
v_gen[1]=256'b1111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000;
v_gen[2]=256'b1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000011111111111111110000000000000000;
v_gen[3]=256'b1111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000;
v_gen[4]=256'b1111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000;
v_gen[5]=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
v_gen[6]=256'b1010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010;
v_gen[7]=256'b1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000;
v_gen[8]=256'b1111111100000000111111110000000000000000000000000000000000000000111111110000000011111111000000000000000000000000000000000000000011111111000000001111111100000000000000000000000000000000000000001111111100000000111111110000000000000000000000000000000000000000;
v_gen[9]=256'b1111000011110000111100001111000000000000000000000000000000000000111100001111000011110000111100000000000000000000000000000000000011110000111100001111000011110000000000000000000000000000000000001111000011110000111100001111000000000000000000000000000000000000;
v_gen[10]=256'b1100110011001100110011001100110000000000000000000000000000000000110011001100110011001100110011000000000000000000000000000000000011001100110011001100110011001100000000000000000000000000000000001100110011001100110011001100110000000000000000000000000000000000;
v_gen[11]=256'b1010101010101010101010101010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000001010101010101010101010101010101000000000000000000000000000000000;
v_gen[12]=256'b1111111100000000000000000000000011111111000000000000000000000000111111110000000000000000000000001111111100000000000000000000000011111111000000000000000000000000111111110000000000000000000000001111111100000000000000000000000011111111000000000000000000000000;
v_gen[13]=256'b1111000011110000000000000000000011110000111100000000000000000000111100001111000000000000000000001111000011110000000000000000000011110000111100000000000000000000111100001111000000000000000000001111000011110000000000000000000011110000111100000000000000000000;
v_gen[14]=256'b1100110011001100000000000000000011001100110011000000000000000000110011001100110000000000000000001100110011001100000000000000000011001100110011000000000000000000110011001100110000000000000000001100110011001100000000000000000011001100110011000000000000000000;
v_gen[15]=256'b1010101010101010000000000000000010101010101010100000000000000000101010101010101000000000000000001010101010101010000000000000000010101010101010100000000000000000101010101010101000000000000000001010101010101010000000000000000010101010101010100000000000000000;
v_gen[16]=256'b1111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000;
v_gen[17]=256'b1100110000000000110011000000000011001100000000001100110000000000110011000000000011001100000000001100110000000000110011000000000011001100000000001100110000000000110011000000000011001100000000001100110000000000110011000000000011001100000000001100110000000000;
v_gen[18]=256'b1010101000000000101010100000000010101010000000001010101000000000101010100000000010101010000000001010101000000000101010100000000010101010000000001010101000000000101010100000000010101010000000001010101000000000101010100000000010101010000000001010101000000000;
v_gen[19]=256'b1100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000;
v_gen[20]=256'b1010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000;
v_gen[21]=256'b1000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000;
v_gen[22]=256'b1111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000;
v_gen[23]=256'b1111000011110000000000000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000011110000111100000000000000000000000000000000000000000000000000001111000011110000000000000000000000000000000000000000000000000000;
v_gen[24]=256'b1100110011001100000000000000000000000000000000000000000000000000110011001100110000000000000000000000000000000000000000000000000011001100110011000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000000000000000000000;
v_gen[25]=256'b1010101010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000;
v_gen[26]=256'b1111000000000000111100000000000000000000000000000000000000000000111100000000000011110000000000000000000000000000000000000000000011110000000000001111000000000000000000000000000000000000000000001111000000000000111100000000000000000000000000000000000000000000;
v_gen[27]=256'b1100110000000000110011000000000000000000000000000000000000000000110011000000000011001100000000000000000000000000000000000000000011001100000000001100110000000000000000000000000000000000000000001100110000000000110011000000000000000000000000000000000000000000;
v_gen[28]=256'b1010101000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000;
v_gen[29]=256'b1100000011000000110000001100000000000000000000000000000000000000110000001100000011000000110000000000000000000000000000000000000011000000110000001100000011000000000000000000000000000000000000001100000011000000110000001100000000000000000000000000000000000000;
v_gen[30]=256'b1010000010100000101000001010000000000000000000000000000000000000101000001010000010100000101000000000000000000000000000000000000010100000101000001010000010100000000000000000000000000000000000001010000010100000101000001010000000000000000000000000000000000000;
v_gen[31]=256'b1000100010001000100010001000100000000000000000000000000000000000100010001000100010001000100010000000000000000000000000000000000010001000100010001000100010001000000000000000000000000000000000001000100010001000100010001000100000000000000000000000000000000000;
v_gen[32]=256'b1111000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000001111000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000001111000000000000000000000000000011110000000000000000000000000000;
v_gen[33]=256'b1100110000000000000000000000000011001100000000000000000000000000110011000000000000000000000000001100110000000000000000000000000011001100000000000000000000000000110011000000000000000000000000001100110000000000000000000000000011001100000000000000000000000000;
v_gen[34]=256'b1010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000;
v_gen[35]=256'b1100000011000000000000000000000011000000110000000000000000000000110000001100000000000000000000001100000011000000000000000000000011000000110000000000000000000000110000001100000000000000000000001100000011000000000000000000000011000000110000000000000000000000;
v_gen[36]=256'b1010000010100000000000000000000010100000101000000000000000000000101000001010000000000000000000001010000010100000000000000000000010100000101000000000000000000000101000001010000000000000000000001010000010100000000000000000000010100000101000000000000000000000;
v_gen[37]=256'b1000100010001000000000000000000010001000100010000000000000000000100010001000100000000000000000001000100010001000000000000000000010001000100010000000000000000000100010001000100000000000000000001000100010001000000000000000000010001000100010000000000000000000;
v_gen[38]=256'b1100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000;
v_gen[39]=256'b1010000000000000101000000000000010100000000000001010000000000000101000000000000010100000000000001010000000000000101000000000000010100000000000001010000000000000101000000000000010100000000000001010000000000000101000000000000010100000000000001010000000000000;
v_gen[40]=256'b1000100000000000100010000000000010001000000000001000100000000000100010000000000010001000000000001000100000000000100010000000000010001000000000001000100000000000100010000000000010001000000000001000100000000000100010000000000010001000000000001000100000000000;
v_gen[41]=256'b1000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000;
v_gen[42]=256'b1111000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000;
v_gen[43]=256'b1100110000000000000000000000000000000000000000000000000000000000110011000000000000000000000000000000000000000000000000000000000011001100000000000000000000000000000000000000000000000000000000001100110000000000000000000000000000000000000000000000000000000000;
v_gen[44]=256'b1010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000;
v_gen[45]=256'b1100000011000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000000000000011000000110000000000000000000000000000000000000000000000000000001100000011000000000000000000000000000000000000000000000000000000;
v_gen[46]=256'b1010000010100000000000000000000000000000000000000000000000000000101000001010000000000000000000000000000000000000000000000000000010100000101000000000000000000000000000000000000000000000000000001010000010100000000000000000000000000000000000000000000000000000;
v_gen[47]=256'b1000100010001000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000000000000000000000;
v_gen[48]=256'b1100000000000000110000000000000000000000000000000000000000000000110000000000000011000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000000001100000000000000110000000000000000000000000000000000000000000000;
v_gen[49]=256'b1010000000000000101000000000000000000000000000000000000000000000101000000000000010100000000000000000000000000000000000000000000010100000000000001010000000000000000000000000000000000000000000001010000000000000101000000000000000000000000000000000000000000000;
v_gen[50]=256'b1000100000000000100010000000000000000000000000000000000000000000100010000000000010001000000000000000000000000000000000000000000010001000000000001000100000000000000000000000000000000000000000001000100000000000100010000000000000000000000000000000000000000000;
v_gen[51]=256'b1000000010000000100000001000000000000000000000000000000000000000100000001000000010000000100000000000000000000000000000000000000010000000100000001000000010000000000000000000000000000000000000001000000010000000100000001000000000000000000000000000000000000000;
v_gen[52]=256'b1100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000011000000000000000000000000000000;
v_gen[53]=256'b1010000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000010100000000000000000000000000000;
v_gen[54]=256'b1000100000000000000000000000000010001000000000000000000000000000100010000000000000000000000000001000100000000000000000000000000010001000000000000000000000000000100010000000000000000000000000001000100000000000000000000000000010001000000000000000000000000000;
v_gen[55]=256'b1000000010000000000000000000000010000000100000000000000000000000100000001000000000000000000000001000000010000000000000000000000010000000100000000000000000000000100000001000000000000000000000001000000010000000000000000000000010000000100000000000000000000000;
v_gen[56]=256'b1000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000;
v_gen[57]=256'b1100000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000;
v_gen[58]=256'b1010000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000;
v_gen[59]=256'b1000100000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000;
v_gen[60]=256'b1000000010000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000;
v_gen[61]=256'b1000000000000000100000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000;
v_gen[62]=256'b1000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000;
v_gen[63]=256'b1000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;
v_gen[64]=256'b1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000;
v_gen[65]=256'b1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[66]=256'b1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[67]=256'b1111111100000000111111110000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000111111110000000011111111000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[68]=256'b1111000011110000111100001111000011110000111100001111000011110000000000000000000000000000000000000000000000000000000000000000000011110000111100001111000011110000111100001111000011110000111100000000000000000000000000000000000000000000000000000000000000000000;
v_gen[69]=256'b1100110011001100110011001100110011001100110011001100110011001100000000000000000000000000000000000000000000000000000000000000000011001100110011001100110011001100110011001100110011001100110011000000000000000000000000000000000000000000000000000000000000000000;
v_gen[70]=256'b1010101010101010101010101010101010101010101010101010101010101010000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010100000000000000000000000000000000000000000000000000000000000000000;
v_gen[71]=256'b1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[72]=256'b1111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[73]=256'b1111000011110000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000111100001111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[74]=256'b1100110011001100110011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011001100110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[75]=256'b1010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[76]=256'b1111111100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[77]=256'b1111000011110000000000000000000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000111100000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[78]=256'b1100110011001100000000000000000011001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000110011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[79]=256'b1010101010101010000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[80]=256'b1111000000000000111100000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[81]=256'b1100110000000000110011000000000011001100000000001100110000000000000000000000000000000000000000000000000000000000000000000000000011001100000000001100110000000000110011000000000011001100000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[82]=256'b1010101000000000101010100000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[83]=256'b1100000011000000110000001100000011000000110000001100000011000000000000000000000000000000000000000000000000000000000000000000000011000000110000001100000011000000110000001100000011000000110000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[84]=256'b1010000010100000101000001010000010100000101000001010000010100000000000000000000000000000000000000000000000000000000000000000000010100000101000001010000010100000101000001010000010100000101000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[85]=256'b1000100010001000100010001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000010001000100010001000100010001000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000;
v_gen[86]=256'b1111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[87]=256'b1111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[88]=256'b1100110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[89]=256'b1010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[90]=256'b1111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[91]=256'b1100110000000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000000001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[92]=256'b1010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[93]=256'b1100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000110000001100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[94]=256'b1010000010100000101000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[95]=256'b1000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[96]=256'b1111000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[97]=256'b1100110000000000000000000000000011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000000000000000000000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[98]=256'b1010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[99]=256'b1100000011000000000000000000000011000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000110000000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[100]=256'b1010000010100000000000000000000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101000000000000000000000101000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[101]=256'b1000100010001000000000000000000010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[102]=256'b1100000000000000110000000000000011000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000001100000000000000110000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[103]=256'b1010000000000000101000000000000010100000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000001010000000000000101000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[104]=256'b1000100000000000100010000000000010001000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000100000000000100010000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[105]=256'b1000000010000000100000001000000010000000100000001000000010000000000000000000000000000000000000000000000000000000000000000000000010000000100000001000000010000000100000001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[106]=256'b1111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[107]=256'b1100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[108]=256'b1010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[109]=256'b1100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[110]=256'b1010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[111]=256'b1000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[112]=256'b1100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[113]=256'b1010000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[114]=256'b1000100000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[115]=256'b1000000010000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[116]=256'b1100000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[117]=256'b1010000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[118]=256'b1000100000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[119]=256'b1000000010000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[120]=256'b1000000000000000100000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[121]=256'b1100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[122]=256'b1010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[123]=256'b1000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[124]=256'b1000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[125]=256'b1000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[126]=256'b1000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[127]=256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[128]=256'b1111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[129]=256'b1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[130]=256'b1111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[131]=256'b1111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[132]=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[133]=256'b1010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[134]=256'b1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[135]=256'b1111111100000000111111110000000000000000000000000000000000000000111111110000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[136]=256'b1111000011110000111100001111000000000000000000000000000000000000111100001111000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[137]=256'b1100110011001100110011001100110000000000000000000000000000000000110011001100110011001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[138]=256'b1010101010101010101010101010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[139]=256'b1111111100000000000000000000000011111111000000000000000000000000111111110000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[140]=256'b1111000011110000000000000000000011110000111100000000000000000000111100001111000000000000000000001111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[141]=256'b1100110011001100000000000000000011001100110011000000000000000000110011001100110000000000000000001100110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[142]=256'b1010101010101010000000000000000010101010101010100000000000000000101010101010101000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[143]=256'b1111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[144]=256'b1100110000000000110011000000000011001100000000001100110000000000110011000000000011001100000000001100110000000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[145]=256'b1010101000000000101010100000000010101010000000001010101000000000101010100000000010101010000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[146]=256'b1100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[147]=256'b1010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000010100000101000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[148]=256'b1000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[149]=256'b1111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[150]=256'b1111000011110000000000000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[151]=256'b1100110011001100000000000000000000000000000000000000000000000000110011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[152]=256'b1010101010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[153]=256'b1111000000000000111100000000000000000000000000000000000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[154]=256'b1100110000000000110011000000000000000000000000000000000000000000110011000000000011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[155]=256'b1010101000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[156]=256'b1100000011000000110000001100000000000000000000000000000000000000110000001100000011000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[157]=256'b1010000010100000101000001010000000000000000000000000000000000000101000001010000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[158]=256'b1000100010001000100010001000100000000000000000000000000000000000100010001000100010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[159]=256'b1111000000000000000000000000000011110000000000000000000000000000111100000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[160]=256'b1100110000000000000000000000000011001100000000000000000000000000110011000000000000000000000000001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[161]=256'b1010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[162]=256'b1100000011000000000000000000000011000000110000000000000000000000110000001100000000000000000000001100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[163]=256'b1010000010100000000000000000000010100000101000000000000000000000101000001010000000000000000000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[164]=256'b1000100010001000000000000000000010001000100010000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[165]=256'b1100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[166]=256'b1010000000000000101000000000000010100000000000001010000000000000101000000000000010100000000000001010000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[167]=256'b1000100000000000100010000000000010001000000000001000100000000000100010000000000010001000000000001000100000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[168]=256'b1000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[169]=256'b1111000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[170]=256'b1100110000000000000000000000000000000000000000000000000000000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[171]=256'b1010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[172]=256'b1100000011000000000000000000000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[173]=256'b1010000010100000000000000000000000000000000000000000000000000000101000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[174]=256'b1000100010001000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[175]=256'b1100000000000000110000000000000000000000000000000000000000000000110000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[176]=256'b1010000000000000101000000000000000000000000000000000000000000000101000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[177]=256'b1000100000000000100010000000000000000000000000000000000000000000100010000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[178]=256'b1000000010000000100000001000000000000000000000000000000000000000100000001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[179]=256'b1100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[180]=256'b1010000000000000000000000000000010100000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[181]=256'b1000100000000000000000000000000010001000000000000000000000000000100010000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[182]=256'b1000000010000000000000000000000010000000100000000000000000000000100000001000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[183]=256'b1000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[184]=256'b1100000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[185]=256'b1010000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[186]=256'b1000100000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[187]=256'b1000000010000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[188]=256'b1000000000000000100000000000000000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[189]=256'b1000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[190]=256'b1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[191]=256'b1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[192]=256'b1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[193]=256'b1111111100000000111111110000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[194]=256'b1111000011110000111100001111000011110000111100001111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[195]=256'b1100110011001100110011001100110011001100110011001100110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[196]=256'b1010101010101010101010101010101010101010101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[197]=256'b1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[198]=256'b1111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[199]=256'b1111000011110000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[200]=256'b1100110011001100110011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[201]=256'b1010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[202]=256'b1111111100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[203]=256'b1111000011110000000000000000000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[204]=256'b1100110011001100000000000000000011001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[205]=256'b1010101010101010000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[206]=256'b1111000000000000111100000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[207]=256'b1100110000000000110011000000000011001100000000001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[208]=256'b1010101000000000101010100000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[209]=256'b1100000011000000110000001100000011000000110000001100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[210]=256'b1010000010100000101000001010000010100000101000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[211]=256'b1000100010001000100010001000100010001000100010001000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[212]=256'b1111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[213]=256'b1111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[214]=256'b1100110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[215]=256'b1010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[216]=256'b1111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[217]=256'b1100110000000000110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[218]=256'b1010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[219]=256'b1100000011000000110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[220]=256'b1010000010100000101000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[221]=256'b1000100010001000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[222]=256'b1111000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[223]=256'b1100110000000000000000000000000011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[224]=256'b1010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[225]=256'b1100000011000000000000000000000011000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[226]=256'b1010000010100000000000000000000010100000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[227]=256'b1000100010001000000000000000000010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[228]=256'b1100000000000000110000000000000011000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[229]=256'b1010000000000000101000000000000010100000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[230]=256'b1000100000000000100010000000000010001000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[231]=256'b1000000010000000100000001000000010000000100000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[232]=256'b1111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[233]=256'b1100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[234]=256'b1010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[235]=256'b1100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[236]=256'b1010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[237]=256'b1000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[238]=256'b1100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[239]=256'b1010000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[240]=256'b1000100000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[241]=256'b1000000010000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[242]=256'b1100000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[243]=256'b1010000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[244]=256'b1000100000000000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[245]=256'b1000000010000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
v_gen[246]=256'b1000000000000000100000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	interface Subifc_Enc_In subifc_in;	
		method Action ma_get_message(Bit#(247) lv_message_in);	
			//(*doc = "note: "fn_mul" is called which will store the returned value into "lv_codeword". " *)
			let lv_codeword = fn_mul(v_gen,lv_message_in);
			
			//(*doc = "fifo:  To store the codeword in FIFO. " *)
			ff_output.enq(lv_codeword);
		endmethod: ma_get_message
	endinterface

	interface Subifc_Enc_Out subifc_out;
		//(*doc = "method: This ActionValue method sends codeword(256 bits) to the channel "*)
		method ActionValue#(Bit#(256)) mav_tx_codeword;
			begin
			//(*doc = "fifo: To remove the contents of the FIFO so that the next set of codeword can be stored. " *)
			ff_output.deq;
			//(*doc = "fifo: To return the contents of FIFO which has the codeword." *)
			return ff_output.first();
			end
		endmethod: mav_tx_codeword
	endinterface
endmodule: mk_rm_encoder

(*synthesize*)
(*doc = "module: Testbench module " *)
module mkTb (Empty);
	//(*doc = "Ifc:  To declare an instance name and instantiate with mk_rm_encoder" *)
	Ifc_rm_encoder ifc_enc<-mk_rm_encoder;
	//(*doc = "note: To declare a vector of 16 elements, each of size 247 bits to store the message before passing into the appropriate method. " *)
	//(*doc = "note:  After 16 cycles, 512 bytes of data will be sent. In the 17 th cycle, 144 bits have to be sent. Append 103 zeroes in order to make it as 247 bits message. Once the codeword for the 17th cycle, take only the bits from the appropriate positions to include the 144 bit message along with the parity bits. " *)
	
	//(*doc = "note: In this code, we are doing it only for two clock cycles.")
	Vector#(2,Bit#(247)) lv_message;
	lv_message[0] = 247'b0000100000010010101101011111111001000001001110001100010010101111001100100010110111000101011100000111100001010111101011011001010110011110011010100110101100110110111110111000011100110100000110011001100000011110001000010001111001010100110100001010100; 
	lv_message[1] = 247'b1000100000010010101101011111111001000001001110001100010010101111001100100010110111000101011100000111100001010111101011011001010110011110011010100110101100110110111110111000011100110100000110011001100000011110001000010001111001010100110100001010100;
			(*doc = "reg: Register to keep track of number of cycles. " *)			
	 		Reg#(Bit#(5)) rg_counter <-mkReg(0);
	
	(*doc = "rule:  To keep sending input message of 247 bits" *)
	rule in (rg_counter<2) ;
			$display($stime," message%d: %b",rg_counter,lv_message[rg_counter]);
			
			//(*doc = "method: The Action method "ma_get_message" is called by passing "lv_message" as argument. " *)
			ifc_enc.subifc_in.ma_get_message(lv_message[rg_counter]);
			//(*doc = "reg: Incrementing the counter to keep track of clock cycles. " *)
			rg_counter <= rg_counter + 1;
	endrule: in
	
	(*doc = "rule: To receive codeword from Encoder" *)
	rule out;
		//(*doc = "method: The ActionValue method "mav_tx_codeword" is called. The returned codeword from the FIFO is stored in "x". " *)
		let lv_x <- ifc_enc.subifc_out.mav_tx_codeword;
		//(*doc = "note: The codeword obtained is displayed. It can be verified if it is a valid codeword by multiplying it with parity check matrix. This can be done in the C program. " *)
		 $display($stime, " codeword: %b ",lv_x);
	endrule: out
	
	(*doc = "rule: To finish simulation " *)
	rule time_finish;	 
		//(*doc = "note: The following code lines are to finish the simulation. " *)
		let lv_time1 <- $stime;
		if(lv_time1 >30)	
			$finish(0);			
	endrule: time_finish		
endmodule: mkTb
endpackage: rm_encoder
